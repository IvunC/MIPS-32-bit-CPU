library ieee; use ieee.std_logic_1164.all; use ieee.numeric_std.all;
--Created By Ivan Contreras
--This File is left as an assignment for the reader.
--JK, since this design was an assignment, I left out the CPU as it is the most vital part
